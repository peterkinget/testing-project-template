* NGSPICE file created from ota_5t.ext - technology: gf180mcuD

.subckt nfet$1 a_30_660# a_254_0# a_n84_0# a_94_0# a_190_660# VSUBS
X0 a_254_0# a_190_660# a_94_0# VSUBS nfet_03v3 ad=1.83p pd=7.22u as=0.78p ps=3.52u w=3u l=0.28u
X1 a_94_0# a_30_660# a_n84_0# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=1.83p ps=7.22u w=3u l=0.28u
.ends

.subckt unit_nmos nfet$1_0/a_30_660# m2_n266_330# m1_n400_n100# m1_300_n100# a_163_0#
+ nfet$1_0/VSUBS
Xnfet$1_0 nfet$1_0/a_30_660# nfet$1_0/VSUBS nfet$1_0/VSUBS m2_n266_330# nfet$1_0/a_30_660#
+ nfet$1_0/VSUBS nfet$1
.ends

.subckt pfet a_254_0# w_n180_n88# a_188_660# a_28_660# a_n92_0# a_94_0#
X0 a_254_0# a_188_660# a_94_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.28u
X1 a_94_0# a_28_660# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.28u
.ends

.subckt unit_pmos m1_311_n100# m2_n264_50# pfet_0/a_28_660# m2_n264_330# m1_n389_n100#
Xpfet_0 m2_n264_50# m2_n264_50# pfet_0/a_28_660# pfet_0/a_28_660# m2_n264_50# m2_n264_330#
+ pfet
.ends

.subckt ota_5t vdd vss i_bias in_n in_p out
Xunit_nmos_0[0|0] i_bias i_bias vss vss vss vss unit_nmos
Xunit_nmos_0[1|0] vss vss vss vss vss vss unit_nmos
Xunit_nmos_0[0|1] i_bias vss vss vss vss vss unit_nmos
Xunit_nmos_0[1|1] in_p m3_n614_1230# vss vss vss vss unit_nmos
Xunit_nmos_0[0|2] i_bias vss vss vss vss vss unit_nmos
Xunit_nmos_0[1|2] in_n out vss vss vss vss unit_nmos
Xunit_nmos_0[0|3] vss vss vss vss unit_nmos_0[0|3]/a_163_0# vss unit_nmos
Xunit_nmos_0[1|3] vss vss vss vss unit_nmos_0[1|3]/a_163_0# vss unit_nmos
Xunit_pmos_0[0|0] vdd vdd vdd vdd vdd unit_pmos
Xunit_pmos_0[1|0] vdd vdd m3_n614_1230# out vdd unit_pmos
Xunit_pmos_0[0|1] vdd vdd m3_n614_1230# out vdd unit_pmos
Xunit_pmos_0[1|1] vdd vdd m3_n614_1230# out vdd unit_pmos
Xunit_pmos_0[0|2] vdd vdd m3_n614_1230# m3_n614_1230# vdd unit_pmos
Xunit_pmos_0[1|2] vdd vdd m3_n614_1230# m3_n614_1230# vdd unit_pmos
Xunit_pmos_0[0|3] vdd vdd vdd vdd vdd unit_pmos
Xunit_pmos_0[1|3] vdd vdd m3_n614_1230# m3_n614_1230# vdd unit_pmos
.ends

